`define module_name i2c_master_driver
