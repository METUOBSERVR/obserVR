module i2c (
    input   A,
    output  B
);
assign  B = A;
endmodule 